module traffic_light (
	input	clk, rst,
	input	ta, tb,
	output	la, lb
);

logic[1:0]	state, nextstate, sb



